`timescale 1ns / 1ps

module VGA_Decoder (
    input  logic       clk,
    input  logic       reset,
    output logic       pclk,
    output logic       h_sync,
    output logic       v_sync,
    output logic [9:0] x_pixel,
    output logic [9:0] y_pixel,
    output logic       DE
);

    //logic pclk;
    logic [9:0] h_counter;
    logic [9:0] v_counter;

    pixel_clk_gen U_P_CLK (.*);

    pixel_counter U_P_COUNTER (.*);

    vga_decoder U_VGA_Decoder (.*);

endmodule     


module pixel_clk_gen (
    input  logic clk,
    input  logic reset,
    output logic pclk
);

    logic [1:0] p_counter;  // 100Mhz => 25Mhz  (/4)

    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            p_counter <= 0;
        end else begin
            if (p_counter == 3) begin
                p_counter <= 0;
                pclk <= 1'b1;
            end else begin
                p_counter <= p_counter + 1;
                pclk <= 1'b0;
            end
        end
    end

endmodule


module pixel_counter (
    input logic pclk,
    input logic reset,
    output logic [9:0] v_counter,
    output logic [9:0] h_counter
);

    localparam H_MAX = 800, V_MAX = 525;  // VGA Spec

    always_ff @(negedge pclk, posedge reset) begin  // horizontal       // negedge에서 처리
        if (reset) begin
            h_counter <= 0;
        end else begin
            if (h_counter == H_MAX - 1) begin
                h_counter <= 0;
            end else begin
                h_counter <= h_counter + 1;
            end
        end
    end

    always_ff @(negedge pclk, posedge reset) begin  // vertical       // negedge에서 처리
        if (reset) begin
            v_counter <= 0;
        end else begin
            if (h_counter == H_MAX - 1) begin
                if (v_counter == V_MAX - 1) begin
                    v_counter <= 0;
                end else begin
                    v_counter <= v_counter + 1;
                end
            end
        end
    end

endmodule


module vga_decoder (
    input  logic pclk,
    input  logic [9:0] h_counter,
    input  logic [9:0] v_counter,
    output logic       h_sync,
    output logic       v_sync,
    output logic [9:0] x_pixel,
    output logic [9:0] y_pixel,
    output logic       DE
);

    localparam H_Display_area = 640;
    localparam H_Front_porch = 16;
    localparam H_Sync_pulse = 96;
    localparam H_Back_porch = 48;
    localparam H_Whole_line = 800;

    localparam V_Display_area = 480;
    localparam V_Front_porch = 10;   
    localparam V_Sync_pulse = 2;
    localparam V_Back_porch = 33;
    localparam V_Whole_frame = 525;

    always_ff @(posedge pclk) begin
        h_sync <= !( (h_counter >= (H_Display_area + H_Front_porch)) && (h_counter < (H_Display_area + H_Front_porch + H_Sync_pulse)) );
        v_sync <= !( (v_counter >= (V_Display_area + V_Front_porch)) && (v_counter < (V_Display_area + V_Front_porch + V_Sync_pulse)) );
        DE <= (h_counter < H_Display_area) && (v_counter < V_Display_area);
        x_pixel <= h_counter;
        y_pixel <= (v_counter >= 525 - 2) ? (v_counter + 2 - 525) : v_counter + 2;
    end
/*   
    assign h_sync = !( (h_counter >= (H_Display_area + H_Front_porch)) && (h_counter < (H_Display_area + H_Front_porch + H_Sync_pulse)) );
    assign v_sync = !( (v_counter >= (V_Display_area + V_Front_porch)) && (v_counter < (V_Display_area + V_Front_porch + V_Sync_pulse)) );

    assign DE = (h_counter < H_Display_area) && (v_counter < V_Display_area);

    assign x_pixel = h_counter;
    assign y_pixel = v_counter;
*/
endmodule
